`timescale 1ns/1ns

module ADD(
    input [31:0]EADD,
    input Ecuatro,
    output reg[31:0]SADD  
);
