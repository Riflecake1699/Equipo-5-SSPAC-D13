`timescale 1ns/1ns
 
 module TB_DATAPATH();

 reg [31:0];
 wire [31:0];

 